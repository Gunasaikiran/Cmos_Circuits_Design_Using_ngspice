***Logic3
.subckt  pass_and 1 2 3 4
.model nmod nmos level=54 version=4.7
M1 1 2 4 4 nmod w=100u l=10u
M2 2 3 4 4 nmod w=100u l=10u
.ends
.subckt  pass_or 1 2 3 4
.model nmod nmos level=54 version=4.7
M1 2 2 4 4 nmod w=100u l=10u
M2 1 3 4 4 nmod w=100u l=10u
.ends
.subckt  invertor 1 2 3
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
M1 3 1 2 2 pmod w=100u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.ends
va 11 0 dc 0v
vb 12 0 dc 0v
vc 13 0 dc 5v
vd 14 0 pulse(0 5 0 0 0 10m 20m)
ve 15 0 dc 0v
vdd 2 0 dc 5v
xb 12 2 16 invertor
xc 13 2 20 invertor
xd 14 2 18 invertor
xcde 21 2 22 invertor
xandb 11 12 16 17 pass_and
xdore 15 14 18 19 pass_or
xdoreandc 19 13 20 21 pass_and
xdoreandcoraandb 17 21 22 23 pass_or
.tran 0.1m 100m
.control
run
set color0 = white
set color1 = black
set xbrushwidth =4.5
plot V(23)
plot V(14)
.endc
.end


