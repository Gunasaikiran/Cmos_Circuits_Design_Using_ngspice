***Trans Analysis
Vin 1 0 pulse(0 5 0 0 0 100ms 200ms)
R1 1 2 6K
C1 2 0 18uF 
.tran 0.2ms 1000ms
.measure tran rtime TRIG V(1) val = 0.5 RISE = 1 TARG V(1) val = 4.5 RISE = 1
.control
run
plot V(1) V(2)
.endc
.end