***DC Analysis
Vin 1 0 5.0V
R1 1 2 8K
R2 2 0 2K 
.dc Vin 0.0 5.0 0.2
.control
run
plot V(1) V(2)
.endc
.end