***DC Analysis
Vin 1 0 5.0V
R1 1 2 1.2K
C1 2 0 0.1uF
L1 2 0 100mH 
.dc Vin 0.0 5.0 0.1
.control
run
plot V(1) V(2)
.endc
.end