*** CMOS INVERTER
Vd 2 0 dc 5V
Vg 1 0 dc 0V
.model nmod nmos level=54 version 4.7
.model pmod pmos level=54 version 4.7
M1 3 1 2 2 pmod w=400u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.dc Vg 0 5 0.1
.control
run
plot V(3) V(1)
.endc
.end

