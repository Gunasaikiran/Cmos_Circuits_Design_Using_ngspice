***AC Analysis
Vin 1 0 dc 0 ac 5V
R1 1 2 6K
C1 2 0 18uF 
.ac dec 10 1 10k
.control
run
plot V(1) V(2)
.endc
.end