***AC Analysis
Vin 1 0 dc 0 ac 5
R1 1 2 8K
R2 2 0 2K 
.ac dec 10 1 10K
.control
run
plot V(1) V(2)
.endc
.end