***Logic1
.subckt  pass_and 1 2 3 4
.model nmod nmos level=54 version=4.7
M1 1 2 4 4 nmod w=100u l=10u
M2 2 3 4 4 nmod w=100u l=10u
.ends
.subckt  pass_or 1 2 3 4
.model nmod nmos level=54 version=4.7
M1 2 2 4 4 nmod w=100u l=10u
M2 1 3 4 4 nmod w=100u l=10u
.ends
.subckt  invertor 1 2 3
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
M1 3 1 2 2 pmod w=100u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.ends
va 11 0 dc 0v
vb 12 0 dc 0v
vc 13 0 dc 0v
vd 14 0 pulse(0 5 0 0 0 10m 20m)
vdd 2 0 dc 5v
xb 12 2 15 invertor
xc 13 2 17 invertor
xd 14 2 19 invertor
xandb 11 12 15 16 pass_and
xabandc 16 13 17 18 pass_and
xabcord 18 14 19 20 pass_or
.tran 0.1m 100m
.control
run
set color0 = white
set color1 = black
set xbrushwidth =4.5
plot V(20)
plot V(14)
.endc
.end


