*** CMOS INVERTER
Vd 2 0 dc 5V
Vg 1 0 pulse(0 5 0 0 0 10m 20m)
.model nmod nmos level=54 version 4.7
.model pmod pmos level=54 version 4.7
M1 3 1 2 2 pmod w=100u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.tran 0.1m 100m
.control
run
plot V(3) V(1)
.endc
.end

