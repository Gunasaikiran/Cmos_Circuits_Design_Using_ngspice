***PMOS CHARACTERSTICS
Vg 1 0 dc -2
Vd 3 0 dc -2.5
V1 3 2 dc 0
.model pmod pmos level=54 version=4.7
M1 0 1 2 2 pmod w=100u 10u
.dc Vg 0 -2.5 -0.1 
.control
run
plot i(V1) xlabel 'Vg' ylabel 'id' 'title' 'transfer character of pmos'
.endc
.end