***Logic2(y=(AB+C(D+E))')
v1 2 0 pulse(0 5 0 0 0 10m 20m)
v2 1 0 dc 5v
v3 3 0 dc 0v
v4 4 0 dc 5v
v5 5 0 dc 5v
vd 11 0 dc 5v
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
m1n 8 2 6 6 nmod w=100u l=10u
m2n 6 1 0 0 nmod w=100u l=10u
m3n 8 3 7 7 nmod w=100u l=10u
m4n 7 4 0 0 nmod w=100u l=10u
m5n 7 5 0 0 nmod w=100u l=10u
m1p 8 3 10 10 pmod w=100u l=10u
m2p 8 5 9 9 pmod w=100u l=10u
m3p 9 4 10 10 pmod w=100u l=10u
m4p 10 2 11 11 pmod w=100u l=10u
m5p 10 1 11 11 pmod w=100u l=10u
.tran 0.1m 100m
.control
run
plot v(8) v(2)
.endc
.end
